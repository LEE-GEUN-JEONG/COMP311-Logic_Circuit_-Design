----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    00:24:17 07/08/2019 
-- Design Name: 
-- Module Name:    test_ex2_mod - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity test_ex2_mod is
	port(a,b : in std_logic;
			y : out std_logic);
end test_ex2_mod;

architecture Behavioral of test_ex2_mod is

begin
	process (a,b)
		begin
		if ( (a='1') and (b='0') ) then
			y <= '1';
			elsif ( (a='0') and (b='1') ) then
			y <= '1';
			else
			y <= '0';
		end if;
	end process;

end Behavioral;

